module filelog